module basicCounter (A,B);

   input A;
   input B;

   assign B=A;

   endmodule
